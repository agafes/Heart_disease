��     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.2�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK
��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR��ExerciseAngina��Oldpeak�et�b�n_features_in_�K
�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h2�f8�����R�(KhNNNNJ����J����K t�b�C              �?�t�bhRh&�scalar���hMC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���K
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hK�
node_count�K��nodes�h(h+K ��h-��R�(KK���h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h~h2�i8�����R�(KhNNNNJ����J����K t�bK ��hh�K��h�h�K��h�h^K��h�h^K ��h�h�K(��h�h^K0��uK8KKt�b�Bx6         ~       	          ����?j8je3�?�           ��@       !                    _@dP,k|��?�            �v@                           �?�H�a��?8            @U@                           �?D^��#��?            �D@                          �]@f���M�?             ?@                          �f@����X�?             @������������������������       �                      @������������������������       �                     @	                          �l@      �?             8@
                          �k@      �?             0@                           �E@�θ�?             *@������������������������       �                     �?                            J@r�q��?
             (@������������������������       �                     @                           �L@����X�?             @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @                           @G@z�G�z�?             $@������������������������       �                      @������������������������       �                      @                          �k@�Ra����?             F@������������������������       �                     A@                           �?      �?	             $@������������������������       �                      @                           @\@      �?              @                          �n@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @"       #       	          ���ٿTc� �?�            �q@������������������������       �                     @$       c                   pq@�	�3�	�?�            @q@%       ,                   @E@ڢPRM�?�            `j@&       +                    �?�n_Y�K�?	             *@'       *                    �?����X�?             @(       )                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @-       <                   `]@ ���3�?|            �h@.       5                    �?�q�q�?             >@/       4                    o@և���X�?
             ,@0       1                    �?���!pc�?             &@������������������������       �                     @2       3                   Pb@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @6       ;                    \@      �?
             0@7       :                   �a@��S�ۿ?	             .@8       9                   @m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?=       ^                    �?�����?h             e@>       O                    �?��S�ۿ?`            �b@?       N                   �b@�T|n�q�?            �E@@       E                   �_@؇���X�?             E@A       D                   �d@�q�q�?             (@B       C                    �K@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @F       K                   �a@��S�ۿ?             >@G       H                    �? 7���B�?             ;@������������������������       �                     4@I       J                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?L       M                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?P       [                    @ 5x ��?E            �Z@Q       Z                   �l@p� V�?B            �Y@R       U                    �?h㱪��?%            �K@S       T                   �c@؇���X�?             @������������������������       �                     �?������������������������       �                     @V       Y                   �a@@��8��?!             H@W       X                    �L@�}�+r��?             3@������������������������       �                     2@������������������������       �                     �?������������������������       �                     =@������������������������       �                     H@\       ]                   �d@      �?             @������������������������       �                     @������������������������       �                     �?_       b                   0a@�q�q�?             2@`       a                   `a@      �?             (@������������������������       �                     @������������������������       �                     @������������������������       �                     @d       s                    �?�G\�c�?)            @P@e       r                    �?��X��?             <@f       k                   �_@��H�}�?             9@g       h                    �H@�8��8��?             (@������������������������       �                      @i       j                   �^@      �?             @������������������������       �                     �?������������������������       �                     @l       q                   8|@�n_Y�K�?             *@m       n                   �a@���!pc�?             &@������������������������       �                     @o       p                   �v@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @t       }                   �d@���@��?            �B@u       |                   �c@b�h�d.�?            �A@v       {                    �?      �?             0@w       x                   �`@�q�q�?             .@������������������������       �                     @y       z                    �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@������������������������       �                      @       �                   �b@
,UP��?�             w@�       �                    @8EGr��?�            �r@�       �                   {@�0����?�            �q@�       �                    �?4_�����?�            �q@�       �                    �R@@�s��?�            @l@�       �                   `_@�8��!�?�             l@�       �       	          ����?��7�K¨?S            @^@�       �                    �?�8��8��?             B@������������������������       �                      @�       �                   �X@г�wY;�?             A@�       �                   �g@�C��2(�?             &@������������������������       �                      @�       �                   @^@�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@������������������������       �        ;            @U@�       �                   �[@,�T�6�?=             Z@�       �                    �D@8����?             7@������������������������       �                     @�       �                   0b@j���� �?	             1@�       �       	             �?�q�q�?             .@�       �                   �m@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �a@ףp=
�?             $@������������������������       �                      @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    @M@H�!b	�?1            @T@�       �                   ``@ qP��B�?            �E@�       �                   Pl@��S�ۿ?             .@������������������������       �                     &@�       �       	             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     <@�       �                    @N@�˹�m��?             C@�       �                   P`@z�G�z�?             $@������������������������       �                     @�       �                    �?�q�q�?             @�       �       	          ���@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �l@h�����?             <@�       �       	          033@ףp=
�?             $@������������������������       �                     @�       �                   �`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             2@������������������������       �                     �?�       �       	             �?�k�'7��?!            �L@������������������������       �                     �?�       �                    �?�X�C�?              L@�       �                    �?�X����?             6@�       �                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	          `ff�?�d�����?             3@�       �                    [@      �?             $@������������������������       �                     @�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     "@�       �                   �`@�IєX�?             A@������������������������       �                     :@�       �                    �?      �?              @������������������������       �                     @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?և���X�?             ,@������������������������       �                     @�       �                    �?z�G�z�?             $@������������������������       �                     �?�       �                   @_@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �       	             @      �?+             Q@�       �                    �?��H�}�?              I@�       �                    �M@z�G�z�?             .@�       �                    �?և���X�?             @������������������������       �                     �?�       �                   �`@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �       	          ����?b�h�d.�?            �A@�       �       	          `ff�?�q�q�?             "@�       �                   �d@z�G�z�?             @�       �                    d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �d@      �?             @������������������������       �                      @������������������������       �                      @�       �                    @K@ȵHPS!�?             :@������������������������       �        
             0@�       �                   �L@�z�G��?             $@������������������������       �                      @�       �                    �L@      �?              @������������������������       �                     @�       �                   @`@      �?             @�       �       	          033�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   g@�����H�?             2@�       �                    @O@�IєX�?
             1@������������������������       �                     *@�       �                   �c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�t�b�values�h(h+K ��h-��R�(KK�KK��h^�B�       Ps@     �z@     @n@      _@      ;@      M@      6@      3@      4@      &@       @      @       @                      @      2@      @      $@      @      $@      @              �?      $@       @      @              @       @      �?       @               @      �?              @                      @       @               @       @       @                       @      @     �C@              A@      @      @       @              @      @      @       @      @                       @              @     �j@     �P@              @     �j@     �N@      f@      A@      @       @      @       @      @      �?              �?      @                      �?              @     �e@      :@      4@      $@      @       @      @       @              @      @      @      @                      @      @              ,@       @      ,@      �?      �?      �?      �?                      �?      *@                      �?      c@      0@     �a@      $@      B@      @      B@      @       @      @      @      @              @      @              @              <@       @      :@      �?      4@              @      �?      @                      �?       @      �?              �?       @                      �?      Z@      @     @Y@       @     �J@       @      @      �?              �?      @             �G@      �?      2@      �?      2@                      �?      =@              H@              @      �?      @                      �?      (@      @      @      @      @                      @      @              C@      ;@      "@      3@      "@      0@      �?      &@               @      �?      @      �?                      @       @      @       @      @      @              �?      @              @      �?                       @              @      =@       @      =@      @      $@      @      $@      @      @              @      @      @                      @              �?      3@                       @     �P@     �r@     �@@     �p@      ;@     0p@      9@      p@      .@     `j@      ,@     `j@      @     �]@      @     �@@       @              �?     �@@      �?      $@               @      �?       @              �?      �?      �?              �?      �?                      7@             @U@      &@     @W@      @      0@              @      @      $@      @      $@      @      �?      @                      �?      �?      "@               @      �?      �?      �?                      �?       @              @     @S@      �?      E@      �?      ,@              &@      �?      @      �?                      @              <@      @     �A@       @       @              @       @      @      �?      @      �?                      @      �?              �?      ;@      �?      "@              @      �?      @              @      �?                      2@      �?              $@     �G@      �?              "@     �G@      @      .@       @      �?              �?       @              @      ,@      @      @              @      @       @      @                       @              "@       @      @@              :@       @      @              @       @               @      �?       @                      �?      @       @      @               @       @      �?              �?       @      �?                       @      A@      A@      @@      2@      @      (@      @      @      �?               @      @              @       @                       @      =@      @      @      @      @      �?      �?      �?      �?                      �?      @               @       @       @                       @      7@      @      0@              @      @               @      @      �?      @              @      �?      �?      �?      �?                      �?       @               @      0@      �?      0@              *@      �?      @              @      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuMhvh(h+K ��h-��R�(KM��h}�B9         x       	          ����?4�5����?�           ��@       7                   �`@�N2��?�            �w@                          �e@8�A�0��?H            �[@                           `@���N8�?             E@                           �?�S����?             C@                          �T@�+e�X�?             9@                           `R@      �?             8@       	                    �D@؇���X�?             5@������������������������       �                     �?
                          �Z@ףp=
�?             4@������������������������       �                      @                          @_@r�q��?	             (@������������������������       �                     @                           �?      �?              @������������������������       �                     �?                           `@����X�?             @������������������������       �                     �?                           @N@r�q��?             @                          @^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@������������������������       �                     @       (                    �?�������?-             Q@                           �?�X���?             F@������������������������       �                     "@       %                    �?և���X�?            �A@                            �?�㙢�c�?             7@������������������������       �                      @!       $                    �G@�����?             5@"       #                   �`@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        	             0@&       '                    @�8��8��?             (@������������������������       �                     &@������������������������       �                     �?)       ,                   (p@      �?             8@*       +       	          hff�?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?-       2                    �?�q�q�?             (@.       1                   q@r�q��?             @/       0                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @3       6                   Pu@�q�q�?             @4       5                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?8       =                   @E@V��T���?�            �p@9       <                    \@@4և���?
             ,@:       ;                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@>       U                    �?������?�            �o@?       B                    �?X���[�?(            �R@@       A                    �?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?C       H                    �?N1���?"            �N@D       G                   �`@�E��ӭ�?	             2@E       F                   �f@     ��?             0@������������������������       �                     *@������������������������       �                     @������������������������       �                      @I       J                    @D@8�$�>�?            �E@������������������������       �                      @K       P                   ``@z�G�z�?            �A@L       M                    g@�z�G��?             4@������������������������       �                     @N       O                    �?և���X�?             ,@������������������������       �                      @������������������������       �                     @Q       R                     M@��S�ۿ?
             .@������������������������       �                     (@S       T                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?V       w                   @g@L�'��T�?i            @f@W       l                    @L@ >�֕�?h            �e@X       a                    �? ��֛�?W            @b@Y       `                   �a@����ȫ�?2            �T@Z       _                    �?�����H�?             "@[       \                   Pa@؇���X�?             @������������������������       �                     @]       ^                   �\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        +            @R@b       k                   `]@      �?%             P@c       j                   `\@z�G�z�?             $@d       i                   @[@�����H�?             "@e       f                    �F@z�G�z�?             @������������������������       �                     @g       h                   @Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     K@m       n                    �?>���Rp�?             =@������������������������       �                     $@o       r                   Hp@p�ݯ��?             3@p       q                    �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?s       v                   �q@؇���X�?             @t       u                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @y       �                    �?61���r�?�            Pv@z       �                    �?N1���?&            �N@{       �                    �?����X�?            �A@|       }                   �Z@�n_Y�K�?             :@������������������������       �                     @~       �                   �m@\X��t�?             7@       �                   �e@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   `\@�q�q�?
             2@������������������������       �                      @�       �                   �q@      �?	             0@������������������������       �                     @�       �                    �?���Q��?             $@�       �                    b@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?      �?             @������������������������       �                     �?�       �       	          ���@�q�q�?             @�       �                     L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                    �H@ȵHPS!�?             :@�       �                    �?�q�q�?             @������������������������       �                      @�       �       	          033�?      �?             @������������������������       �                      @������������������������       �                      @�       �                    \@P���Q�?             4@�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     2@�       �                    @E@P�0�e��?�            �r@�       �                    �?���Q��?             4@�       �                    �?�8��8��?             (@������������������������       �                     "@�       �                    c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �l@      �?              @������������������������       �                     @�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?�                         pv@�	��X�?�            @q@�       �                   P`@�t�o}�?�            q@�       �       	          `ff@     ��?M             `@�       �                   Ph@����?E            @\@�       �       	          033�?�}�+r��?             C@������������������������       �                     2@�       �                    �?ףp=
�?             4@�       �                    W@؇���X�?	             ,@������������������������       �                     �?�       �                    �?$�q-�?             *@�       �       	              @؇���X�?             @�       �                   `_@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?��n�?+            �R@�       �                   �[@H%u��?             9@�       �                   `n@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   �j@�}�+r��?             3@�       �       	          pff�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             0@�       �                    �?H.�!���?             I@�       �                    �?������?            �B@������������������������       �                     @�       �                   0i@�r����?             >@������������������������       �                      @�       �                   �`@@4և���?             <@������������������������       �                     6@�       �                    �?�q�q�?             @������������������������       �                     @�       �                    @K@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �[@��
ц��?             *@������������������������       �                      @�       �                   �\@���|���?             &@������������������������       �                      @�       �                   �b@�<ݚ�?             "@�       �       	             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       	             
@�q�q�?             .@�       �                    �?�n_Y�K�?             *@�       �                    �?�����H�?             "@�       �                   8p@      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?�������?b             b@�       �                   `b@�t����?             1@������������������������       �                     (@�       �                   �d@���Q��?             @�       �                   `o@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�                          �R@     ��?U             `@�       �       	          ����?��b�h8�?T            �_@�       �                    �?z�G�z�?             9@�       �                    �K@�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                    �?      �?             0@�       �                   ``@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @������������������������       �                     @�                          �c@г�wY;�?F            �Y@�       �       	          ����?p���?D             Y@�       �                   �Q@������?            �D@�       �                     N@r�q��?             (@�       �                   �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     =@������������������������       �        *            �M@                        �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMKK��h^�BP       �t@     y@     p@      ^@     �F@     @P@      $@      @@      @      @@      @      3@      @      2@      @      2@      �?               @      2@               @       @      $@              @       @      @              �?       @      @      �?              �?      @      �?       @      �?                       @              @      @                      �?              *@      @             �A@     �@@      =@      .@      "@              4@      .@      3@      @               @      3@       @      @       @               @      @              0@              �?      &@              &@      �?              @      2@      �?      &@              &@      �?              @      @      �?      @      �?       @               @      �?                      @      @       @      @      �?      @                      �?              �?     �j@     �K@      �?      *@      �?       @      �?                       @              &@     `j@      E@      G@      =@      *@      �?      *@                      �?     �@@      <@      @      *@      @      *@              *@      @               @              <@      .@               @      <@      @      ,@      @      @               @      @       @                      @      ,@      �?      (@               @      �?       @                      �?     �d@      *@     �d@      $@     �a@      @     @T@      �?       @      �?      @      �?      @               @      �?              �?       @               @             @R@              O@       @       @       @       @      �?      @      �?      @              �?      �?      �?                      �?      @                      �?      K@              6@      @      $@              (@      @      &@      �?      &@                      �?      �?      @      �?       @               @      �?                      @              @      S@     �q@     �@@      <@      $@      9@      $@      0@              @      $@      *@      @      �?              �?      @              @      (@       @              @      (@              @      @      @      @      @      @                      @      �?      @              �?      �?       @      �?      �?              �?      �?                      �?              "@      7@      @      @       @       @               @       @               @       @              3@      �?      �?      �?              �?      �?              2@             �E@     �o@       @      (@      �?      &@              "@      �?       @      �?                       @      @      �?      @              @      �?      @                      �?     �A@      n@      @@      n@      5@     �Z@      0@     @X@       @      B@              2@       @      2@       @      (@      �?              �?      (@      �?      @      �?      @              @      �?                       @              @              @      ,@     �N@      @      6@       @      @       @                      @      �?      2@      �?       @      �?                       @              0@      &@     �C@      @     �@@              @      @      :@       @               @      :@              6@       @      @              @       @      �?       @                      �?      @      @               @      @      @               @      @       @      @       @      @                       @      @              @      $@      @       @      �?       @      �?      @               @      �?      �?              �?      �?                      @      @                       @      &@     �`@       @      .@              (@       @      @       @      �?       @                      �?               @      "@     �]@       @     �]@      @      4@      @      @      @                      @       @      ,@       @      &@              &@       @                      @      @     �X@       @     �X@       @     �C@       @      $@       @       @       @                       @               @              =@             �M@      �?      �?      �?                      �?      �?              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK녔h}�Bh3         2                    �?p�Vv���?�           ��@              	          ����?�>�p���?Y             b@                          �Q@�����H�?4            @T@                          a@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?�:�^���?1            �S@                           d@�t����?
             1@	       
                     J@8�Z$���?             *@������������������������       �                      @                           ]@���Q��?             @������������������������       �                      @                           �?�q�q�?             @                          �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                          @d@      �?             @������������������������       �                     @������������������������       �                     �?                           �?�]0��<�?'            �N@������������������������       �        "             J@                           �L@�<ݚ�?             "@                           a@�q�q�?             @                           �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       -                    �?     ��?%             P@       $                    �?������?            �F@        !                   �R@j���� �?             1@������������������������       �                     @"       #       	          `ff@����X�?             ,@������������������������       �                     $@������������������������       �                     @%       ,       	          ����?@4և���?             <@&       '                    �?"pc�
�?             &@������������������������       �                     @(       )                   �m@����X�?             @������������������������       �                     �?*       +                   @_@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     1@.       1       	          ����?�}�+r��?             3@/       0                   `c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@3       �                    �?~�.���?�           h�@4       ?                   �_@|�38���?�            �t@5       6                    �?���J��?C            �Y@������������������������       �        -            @Q@7       8       	          033�?�FVQ&�?            �@@������������������������       �                     9@9       :                   @`@      �?              @������������������������       �                     �?;       >                    �?؇���X�?             @<       =                   `]@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @@       s                    �?P̏����?�            �l@A       T                   �`@�i#[��?9             U@B       O                   �k@8^s]e�?             =@C       F                   �Y@���Q��?             4@D       E                    �?����X�?             @������������������������       �                     @������������������������       �                      @G       L                    �?�θ�?
             *@H       K                   pi@ףp=
�?             $@I       J                   �g@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @M       N                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?P       S                    �G@�����H�?             "@Q       R                   Hy@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @U       l                   �n@N{�T6�?#            �K@V       g                   �e@���y4F�?             C@W       Z                    �D@6YE�t�?            �@@X       Y       	          @33�?�q�q�?             @������������������������       �                     �?������������������������       �                      @[       f                   pk@ףp=
�?             >@\       e       	          hff�?r�q��?
             2@]       d                    �?�t����?	             1@^       c       	          ����?�r����?             .@_       `                   �b@"pc�
�?             &@������������������������       �                     @a       b                   �\@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@h       i                    �D@���Q��?             @������������������������       �                      @j       k                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @m       r                   b@������?             1@n       q                   �z@�q�q�?             @o       p                    @N@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@t       �                   (q@�5?,R�?b             b@u       �                   q@0w-!��?F             Y@v       �                    �?�^'�ë�?E            @X@w       �                   �e@      �?6             T@x       y                   i@���!���?5            �S@������������������������       �                     2@z       �                   @j@f>�cQ�?(            �N@{       |       	             �?����X�?             @������������������������       �                     �?}       �                   �i@r�q��?             @~              	          033�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �       	            �?�>����?#             K@�       �       	          ����?      �?             @�       �                   `a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   �[@`2U0*��?              I@������������������������       �                     ,@�       �                    �J@�X�<ݺ?             B@�       �                    @J@�r����?             .@�       �                   �m@$�q-�?	             *@������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     5@������������������������       �                     �?������������������������       �                     1@������������������������       �                     @������������������������       �                     F@�       �       	          ����?��?�            0p@�       �                    @�}���?x             h@�       �                   �X@,�"���?l            @e@�       �                    @G@���!pc�?	             &@������������������������       �                      @�       �                   @`@�����H�?             "@�       �                   `V@z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �O@���C��?c            �c@�       �                    �?      �?              @������������������������       �                      @�       �                   �`@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �K@tX�}}��?]            �b@�       �                   �g@���#�İ?F            �]@�       �                    @H@ ���J��?E            @]@�       �                    �G@xL��N�?+            �R@�       �                   �a@����e��?&            �P@�       �                   `a@��S�ۿ?	             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �                    �I@�       �                   �d@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                    �E@������������������������       �                     �?�       �                   �a@�q�q�?            �@@�       �       	          ����?�G�z��?             4@�       �                    �?�q�q�?             .@�       �                   �i@X�<ݚ�?             "@������������������������       �                      @�       �                   �a@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    @L@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �P@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@�       �                   �c@�û��|�?             7@�       �                   �p@��.k���?	             1@�       �                   `Q@      �?             (@������������������������       �                     @������������������������       �                     "@������������������������       �                     @������������������������       �                     @�       �                   P`@r�q��?0            �P@�       �                    `@�LQ�1	�?             7@�       �       	          ��� @�d�����?             3@�       �                   �^@�eP*L��?
             &@�       �                   �o@����X�?             @�       �                   �\@      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �Z@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �       	             @      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     E@Du9iH��?            �E@������������������������       �                     �?�       �                   pb@���N8�?             E@������������������������       �                    �@@�       �                   �h@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h^�B�       @t@     �y@     �Y@     �E@      R@      "@      �?       @      �?                       @     �Q@      @      (@      @      &@       @       @              @       @       @              �?       @      �?      �?              �?      �?                      �?      �?      @              @      �?             �M@       @      J@              @       @      @       @      @      �?      @                      �?              �?      @              >@      A@      (@     �@@      $@      @              @      $@      @      $@                      @       @      :@       @      "@              @       @      @      �?              �?      @      �?                      @              1@      2@      �?      @      �?      @                      �?      .@             �k@     �v@      M@      q@       @      Y@             @Q@       @      ?@              9@       @      @      �?              �?      @      �?      @              @      �?                      @      L@     �e@     �E@     �D@      "@      4@       @      (@      @       @      @                       @      @      $@      �?      "@      �?      �?              �?      �?                       @       @      �?       @                      �?      �?       @      �?       @      �?                       @              @      A@      5@      >@       @      <@      @      �?       @      �?                       @      ;@      @      .@      @      .@       @      *@       @      "@       @      @              @       @      @                       @      @               @                      �?      (@               @      @               @       @      �?              �?       @              @      *@      @       @      @      �?      @                      �?              �?              &@      *@     ``@      *@     �U@      $@     �U@      $@     �Q@      "@     �Q@              2@      "@      J@      @       @              �?      @      �?      @      �?      @                      �?       @              @      I@       @       @      �?       @               @      �?              �?               @      H@              ,@       @      A@       @      *@      �?      (@               @      �?      @              @      �?              �?      �?              �?      �?                      5@      �?                      1@      @                      F@     �d@     �W@      c@      D@      b@      :@      @       @       @              �?       @      �?      @      �?      �?      �?                      �?              @              @     �a@      2@      @      @       @              @      @              @      @              a@      .@     �\@      @     �\@      @     �Q@      @     @P@      �?      ,@      �?      ,@                      �?     �I@              @       @      @                       @     �E@                      �?      6@      &@      "@      &@      @      $@      @      @               @      @      @      @                      @      �?      @      �?                      @      @      �?      @                      �?      *@              "@      ,@      "@       @      "@      @              @      "@                      @              @      &@     �K@       @      .@      @      ,@      @      @       @      @       @       @              �?       @      �?      �?              �?      �?              �?      �?                      @      @      �?              �?      @                       @      @      �?       @              �?      �?              �?      �?              @      D@      �?               @      D@             �@@       @      @       @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK���h}�Bx6         r                   �`@U�ք�?�           ��@       C                   �`@�~6�]�?�            @u@       "                    �?�G�z��?n             d@                           �?      �?/             Q@                           �?�"U����?%            �I@                          p`@�Q����?             D@                           �?�s��:��?             C@       	       	          ����?��S�ۿ?             .@������������������������       �        	             (@
                          �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?8����?             7@                           [@$�q-�?             *@                          �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             &@                          �Z@���Q��?             $@������������������������       �                     @                          �Y@؇���X�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     &@                           �?�t����?
             1@������������������������       �                     �?              	          ����?      �?	             0@������������������������       �                     "@        !                    �L@؇���X�?             @������������������������       �                     @������������������������       �                     �?#       B                    `@��A��??             W@$       3                   �^@z���=��?4            @S@%       (                    [@@4և���?             E@&       '       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @)       0                   Hs@�7��?            �C@*       +                    @L@��?^�k�?            �A@������������������������       �                     5@,       /                    \@@4և���?
             ,@-       .                    Y@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@1       2                   �t@      �?             @������������������������       �                     �?������������������������       �                     @4       7                    �?����X�?            �A@5       6                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @8       ?       	          ����?V�a�� �?             =@9       :                   �Y@�n_Y�K�?             *@������������������������       �                     @;       <       	          ����?      �?              @������������������������       �                      @=       >                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?@       A                   @_@      �?	             0@������������������������       �                     �?������������������������       �                     .@������������������������       �                     .@D       M                    �G@4?,R��?k            �f@E       F                   @a@�z�G��?             $@������������������������       �                     �?G       H                    �?�<ݚ�?             "@������������������������       �                     @I       J                    �?      �?             @������������������������       �                     �?K       L                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @N       c       	          033�?�̨�`<�?d            @e@O       b                    �?      �?             F@P       _       	          ����?��>4և�?             <@Q       ^                     O@���!pc�?             6@R       Y                    �?���Q��?
             .@S       T                    �?�����H�?             "@������������������������       �                     @U       X                    �?r�q��?             @V       W                     K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @Z       [                    �?r�q��?             @������������������������       �                     @\       ]                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @`       a                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             0@d       q                    `R@�X�<ݺ?I            �_@e       j                    `@`J����?H            �^@f       g                    @@���a��?C            �\@������������������������       �        A            �[@h       i                    �?      �?             @������������������������       �                     �?������������������������       �                     @k       p                    @N@      �?              @l       m       	          ����?      �?             @������������������������       �                      @n       o       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @s       �                    �?�����?           �x@t       �                    @L@�z�G��?�            �t@u       �       	             @���0��?�            �m@v       �                   @g@B�Y��f�?�            �l@w       �                   �`@&^�r���?�            @l@x       �                   `]@�Z��=��?j            �c@y       z                   pb@      �?             D@������������������������       �                     .@{       |                   0c@���Q��?             9@������������������������       �                     @}       �                   �p@�X����?             6@~                           �?     ��?             0@������������������������       �                     @�       �                   �i@�z�G��?             $@������������������������       �                     @�       �                    �F@      �?             @������������������������       �                      @�       �                    d@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?|�űN�?P            @]@������������������������       �                     F@�       �                    �G@L������?5            @R@�       �                    �?���N8�?             E@������������������������       �                     �?�       �                    @��Y��]�?            �D@������������������������       �                     D@������������������������       �                     �?�       �                    �?�n`���?             ?@�       �                   �^@      �?
             (@�       �                    b@z�G�z�?             @������������������������       �                      @�       �                     I@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    `@����X�?             @������������������������       �                     @�       �       	          433�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     3@�       �                   �`@�G�5��?1            @Q@�       �                   @c@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    @Z���c��?,            �O@�       �                    �?�:�B��?)            �M@������������������������       �                     &@�       �       	          @33�?�q�q�?"             H@�       �                   �f@�C��2(�?            �@@�       �                   xp@`Jj��?             ?@������������������������       �                     2@�       �                    �?8�Z$���?             *@�       �                   �p@�8��8��?
             (@�       �                    @E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?�       �                   g@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?��S���?             .@������������������������       �                      @�       �                    �G@�n_Y�K�?             *@������������������������       �                     @�       �                     J@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @�       �                   `f@      �?             @�       �       	          `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?z�G�z�?	             $@������������������������       �                     �?�       �                   n@�����H�?             "@������������������������       �                     @�       �                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �j@��c:�?7             W@�       �                   @a@     ��?             0@������������������������       �                      @�       �                    @N@      �?              @������������������������       �                     @������������������������       �                     @�       �       	          `ff�?���=A�?+             S@�       �                    �?*O���?             B@�       �       	             �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �q@������?             >@�       �                    �?؇���X�?             5@������������������������       �                     "@�       �                    �M@      �?             (@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?X�<ݚ�?             "@������������������������       �                     @�       �                   0b@�q�q�?             @������������������������       �                      @�       �                   ht@      �?             @������������������������       �                     �?�       �                   u@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?P���Q�?             D@������������������������       �                     >@�       �                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @�       �                    �?     ��?)             P@������������������������       �                     B@�       �                   �o@��X��?             <@�       �                    @z�G�z�?             4@�       �                   �O@�S����?             3@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @M@      �?             0@������������������������       �                     (@�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �q@      �?              @������������������������       �                     @�       �                   c@      �?             @������������������������       �                     �?������������������������       �                     @�t�b�l!     h�h(h+K ��h-��R�(KK�KK��h^�B�        t@     �y@      R@     �p@     �G@     @\@      A@      A@      @@      3@      5@      3@      5@      1@      ,@      �?      (@               @      �?              �?       @              @      0@      �?      (@      �?      �?      �?                      �?              &@      @      @              @      @      �?      �?      �?              �?      �?              @                       @      &@               @      .@      �?              �?      .@              "@      �?      @              @      �?              *@     �S@      *@      P@      @     �C@      �?       @      �?                       @       @     �B@      �?      A@              5@      �?      *@      �?      @              @      �?                      $@      �?      @      �?                      @      $@      9@      @       @               @      @              @      7@      @       @              @      @      @               @      @      �?      @                      �?      �?      .@      �?                      .@              .@      9@     `c@      @      @              �?      @       @      @               @       @              �?       @      �?              �?       @              2@      c@      &@     �@@      &@      1@      @      0@      @      "@      �?       @              @      �?      @      �?       @               @      �?                      @      @      �?      @               @      �?       @                      �?              @      @      �?              �?      @                      0@      @     �]@      @     �]@      �?     �\@             �[@      �?      @      �?                      @      @      @      @      �?       @              �?      �?              �?      �?                      @      @             @o@      b@     �l@     �X@      h@     �F@     �g@     �B@     �g@     �A@     `a@      2@      >@      $@      .@              .@      $@              @      .@      @      "@      @      @              @      @              @      @      @       @              �?      @      �?                      @      @             @[@       @      F@             @P@       @      D@       @              �?      D@      �?      D@                      �?      9@      @      @      @      @      �?       @               @      �?       @                      �?       @      @              @       @      �?       @                      �?      3@              J@      1@       @      @              @       @              I@      *@     �H@      $@      &@              C@      $@      >@      @      =@       @      2@              &@       @      &@      �?      �?      �?      �?                      �?      $@                      �?      �?      �?              �?      �?               @      @               @       @      @      @              @      @              @      @              �?      @      �?      �?              �?      �?                       @               @       @       @      �?              �?       @              @      �?      �?      �?                      �?      C@      K@      *@      @       @              @      @      @                      @      9@     �I@      7@      *@      �?      @              @      �?              6@       @      2@      @      "@              "@      @      �?      @              @      �?               @              @      @              @      @       @       @               @       @      �?              �?       @               @      �?               @      C@              >@       @       @       @                       @      3@     �F@              B@      3@      "@      0@      @      0@      @      �?       @               @      �?              .@      �?      (@              @      �?              �?      @                      �?      @      @              @      @      �?              �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuM	hvh(h+K ��h-��R�(KM	��h}�B�9         �       	          ����?4�5����?�           ��@       7                    @J@�Ff��K�?�            x@                           �?H芦��?�            �j@                          i@J�����?/            @S@                           �?��� ��?             ?@                          �Z@��s����?             5@������������������������       �                      @       	                     H@�KM�]�?
             3@������������������������       �                     .@
                           @I@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     $@                            B@���j��?             G@������������������������       �                     @                          �Z@>��C��?            �E@������������������������       �                     @                          hp@z�G�z�?             D@                          �Y@�>����?             ;@                           l@      �?              @������������������������       �                     �?������������������������       �                     �?                          �b@`2U0*��?             9@������������������������       �                     8@������������������������       �                     �?                          �a@�n_Y�K�?             *@������������������������       �                     @                          0d@r�q��?             @������������������������       �                     @������������������������       �                     �?                            �?���.�6�?W            @a@������������������������       �                    �G@!       .                   `]@�ɮ����?<            �V@"       -                   `\@�q�q�?
             .@#       ,                    �?����X�?	             ,@$       %       	          ������	j*D�?             *@������������������������       �                     �?&       +                   �o@�q�q�?             (@'       *                   @[@�����H�?             "@(       )                    i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?/       0                   `a@�}�+r��?2             S@������������������������       �                     F@1       2                   �b@      �?             @@������������������������       �                     &@3       4                   �d@��s����?             5@������������������������       �                     @5       6                   pe@�X�<ݺ?             2@������������������������       �                     �?������������������������       �                     1@8       o                    �?k�q��?s            @e@9       F                   �a@�������?S             ]@:       C                    �?8����?             7@;       @                   �_@���Q��?             .@<       =                   �`@�����H�?             "@������������������������       �                     @>       ?                    �?      �?              @������������������������       �                     �?������������������������       �                     �?A       B                    @r�q��?             @������������������������       �                     @������������������������       �                     �?D       E                   �`@      �?              @������������������������       �                     @������������������������       �                     �?G       n                   �g@��!���?D            @W@H       O                    �?@S�)�q�?C            �V@I       N                    �?�g�y��?             ?@J       K                   d@�����H�?             "@������������������������       �                     @L       M                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     6@P       m                   xt@������?/             N@Q       ^                    �?>���Rp�?.             M@R       U                   �\@\X��t�?             7@S       T                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?V       ]       	          @33�?�t����?             1@W       X                   �f@�eP*L��?	             &@������������������������       �                      @Y       Z                   @^@X�<ݚ�?             "@������������������������       �                     @[       \                   �n@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @_       d                    b@(N:!���?            �A@`       a       	          pff�?`2U0*��?             9@������������������������       �                     4@b       c                     L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?e       l                   �p@�z�G��?	             $@f       g                    X@�<ݚ�?             "@������������������������       �                     �?h       k                   c@      �?              @i       j                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @p       �                   �b@�{��?��?              K@q       v                    �?8��8���?             H@r       u                   �^@���Q��?             @s       t                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @w       |                   �`@X�EQ]N�?            �E@x       {                   �Z@ ��WV�?             :@y       z                    �O@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@}       �       	             �?������?             1@~       �                    �?؇���X�?	             ,@       �                   �T@����X�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �c@�q�q�?             @������������������������       �                      @�       �                     Q@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �b@�?ʵ���?�            �u@�       �       	          ����?؇���X�?�            �q@�       �                   �`@~X�<��?2             R@�       �                    �E@Z�K�D��?            �G@������������������������       �                      @�       �                    W@��Zy�?            �C@�       �                    `@�����H�?             "@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          `ff�?��S���?             >@������������������������       �                     �?�       �                   @Z@П[;U��?             =@������������������������       �                     @�       �                    �K@��H�}�?             9@�       �                   �`@և���X�?
             ,@�       �                    �?z�G�z�?             $@������������������������       �                     �?�       �                    �?�����H�?             "@�       �                   @_@r�q��?             @�       �                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                     P@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                    �?HP�s��?             9@������������������������       �                     4@�       �                    @L@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?ܾ�z�<�?�             j@�       �                   ``@���`uӽ?k             d@�       �                    �?�y��*�?*             M@�       �                    �?���!pc�?             &@�       �                   �`@���Q��?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       	             @dP-���?#            �G@�       �                    �?P���Q�?             D@�       �                   `_@�8��8��?             8@������������������������       �                     .@�       �                   j@�<ݚ�?             "@�       �       	             @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     0@�       �                   �Z@����X�?             @������������������������       �                     �?�       �                   �_@r�q��?             @�       �                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   P`@ f^8���?A            �Y@�       �                   �r@����ȫ�?1            �T@������������������������       �        '            �O@�       �                    �?�}�+r��?
             3@������������������������       �        	             2@������������������������       �                     �?�       �                   p`@�����?             5@������������������������       �                     �?�       �                   �c@P���Q�?             4@������������������������       �                     0@�       �                    @O@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?��|�5��?            �G@�       �                   �n@؇���X�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   0g@      �?             D@�       �                    @�d�����?             3@�       �                    ]@8�Z$���?	             *@�       �                    �?�q�q�?             @������������������������       �                      @�       �                     O@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   @_@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     5@�             	             @ꮃG��?/            @Q@�       �                    �?N{�T6�?%            �K@�       �                   �g@���"͏�?            �B@������������������������       �                      @�       �                    �?z�G�z�?            �A@������������������������       �                     (@�       �                    �L@8����?             7@�       �                   �q@r�q��?             2@�       �                   �\@���!pc�?	             &@������������������������       �                      @�       �                   �e@�����H�?             "@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   pc@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�                          �?�q�q�?             2@�                           q@$�q-�?	             *@������������������������       �                     &@                        pd@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                         �?@4և���?
             ,@������������������������       �                     &@                        �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KM	KK��h^�B�       �t@     y@      p@     �_@     �d@     �H@     �B@      D@      @      ;@      @      1@       @               @      1@              .@       @       @       @                       @              $@     �@@      *@              @     �@@      $@              @     �@@      @      9@       @      �?      �?              �?      �?              8@      �?      8@                      �?       @      @      @              �?      @              @      �?              `@      "@     �G@             �T@      "@      $@      @      $@      @      "@      @      �?               @      @       @      �?      �?      �?      �?                      �?      @                      @      �?                      �?      R@      @      F@              <@      @      &@              1@      @              @      1@      �?              �?      1@              W@     �S@     @T@     �A@      @      0@      @      "@      �?       @              @      �?      �?              �?      �?              @      �?      @                      �?      �?      @              @      �?             �R@      3@     �R@      1@      >@      �?       @      �?      @               @      �?       @                      �?      6@              F@      0@      F@      ,@      *@      $@      �?      @              @      �?              (@      @      @      @       @              @      @      @              �?      @              @      �?              @              ?@      @      8@      �?      4@              @      �?      @                      �?      @      @      @       @              �?      @      �?      �?      �?      �?                      �?      @                      �?               @               @      &@     �E@      @     �D@       @      @       @      �?       @                      �?               @      @      C@      �?      9@      �?      @              @      �?                      2@      @      *@       @      (@       @      @       @      �?              �?       @                      @              @       @      �?       @                      �?      @       @       @               @       @       @                       @     �R@      q@      D@      n@      3@     �J@      1@      >@               @      1@      6@      �?       @              @      �?       @               @      �?              0@      ,@              �?      0@      *@              @      0@      "@      @       @       @       @      �?              �?       @      �?      @      �?      �?              �?      �?                      @              @      @              $@      �?      $@                      �?       @      7@              4@       @      @       @                      @      5@     `g@      $@     �b@      @     �I@      @       @      @       @      �?       @      �?                       @       @                      @      @     �E@       @      C@       @      6@              .@       @      @       @      �?       @                      �?              @              0@       @      @      �?              �?      @      �?      �?              �?      �?                      @      @      Y@      �?     @T@             �O@      �?      2@              2@      �?               @      3@      �?              �?      3@              0@      �?      @              @      �?              &@      B@      @      �?      @               @      �?       @                      �?      @     �A@      @      ,@       @      &@       @      @               @       @       @               @       @                      @      @      @      @                      @              5@     �A@      A@      A@      5@      <@      "@               @      <@      @      (@              0@      @      .@      @       @      @               @       @      �?      @              �?      �?      �?                      �?      @              �?      @      �?                      @      @      (@      �?      (@              &@      �?      �?      �?                      �?      @              �?      *@              &@      �?       @      �?                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuMhvh(h+K ��h-��R�(KM��h}�B88         �       	          ����?6������?�           ��@                          @E@��_���?�             w@       
                    �?�S����?$            �L@                           �? >�֕�?            �A@������������������������       �                     9@                           [@z�G�z�?             $@������������������������       �                     @       	                   �]@���Q��?             @������������������������       �                      @������������������������       �                     @                          �_@�X����?             6@                          `]@@4և���?             ,@������������������������       �                     "@                           �?z�G�z�?             @������������������������       �                     @                          �^@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?      �?              @������������������������       �                     @������������������������       �                      @       W                   �n@�W�o���?�            ps@       >                    �?\[j��?v             g@       =                    �?��0u���?&             N@       $                   �]@�BbΊ�?$             M@       #                   j@      �?             0@       "                    �?z�G�z�?             $@                           @G@����X�?             @������������������������       �                     @                           �?�q�q�?             @������������������������       �                     �?        !                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @%       :                   �e@r�q��?             E@&       /                   pf@�ݜ�?            �C@'       .                    �?և���X�?             @(       )                    �L@z�G�z�?             @������������������������       �                      @*       -                     O@�q�q�?             @+       ,                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @0       5                   �i@      �?             @@1       4       	          @33�?؇���X�?             @2       3                    �L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @6       7                    @O@`2U0*��?             9@������������������������       �        	             4@8       9                    �O@z�G�z�?             @������������������������       �                     �?������������������������       �                     @;       <                     F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @?       B                   �W@0{�v��?P            @_@@       A                    �?      �?             @������������������������       �                     @������������������������       �                     @C       T                    `P@hx<?v��?N            �]@D       M                   �l@ T���v�?K            @\@E       L                   �a@�q�q�??             X@F       K                   p`@Pa�	�?            �@@G       H                    �?@4և���?             ,@������������������������       �        	             (@I       J                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     3@������������������������       �        )            �O@N       O                    �?�t����?             1@������������������������       �                     &@P       Q                   �l@�q�q�?             @������������������������       �                     �?R       S                    @G@z�G�z�?             @������������������������       �                     @������������������������       �                     �?U       V                    �?      �?             @������������������������       �                     @������������������������       �                     @X       u                    �?X�Cc�?Q            �_@Y       Z                   �Z@�d�����?             C@������������������������       �                     �?[       b                    @F@���"͏�?            �B@\       a                    �D@�C��2(�?             &@]       `                    �?z�G�z�?             @^       _                    _@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @c       j                    �?�	j*D�?             :@d       e                     J@���Q��?             $@������������������������       �                     @f       g                   �b@և���X�?             @������������������������       �                      @h       i                    �?���Q��?             @������������������������       �                      @������������������������       �                     @k       n                   Xp@      �?	             0@l       m                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?o       t                   b@@4և���?             ,@p       s                    @J@z�G�z�?             @q       r                   �p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@v       w                    Z@
�GN��?:             V@������������������������       �                     @x       �                    �K@P�;�&��?8            @U@y       ~                   `]@     ��?(             P@z       {                   �e@���|���?             &@������������������������       �                     @|       }                   p@z�G�z�?             @������������������������       �                     �?������������������������       �                     @       �                    @�&=�w��?#            �J@�       �                    �? pƵHP�?"             J@������������������������       �                     E@�       �                    �?ףp=
�?             $@������������������������       �                     @�       �                    @I@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   �b@�ՙ/�?             5@�       �                   ht@     ��?             0@�       �                   �`@؇���X�?             ,@�       �                    �L@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@�       �                   u@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?xƅd�?�            �v@�       �                    �? �&�T�?�            @q@�       �       	          033�?���Q��?              I@�       �                   @[@      �?             @@������������������������       �                     @�       �                    �?д>��C�?             =@�       �                   �`@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �        	             4@�       �                    �?�q�q�?             2@������������������������       �                     (@������������������������       �                     @�       �                   �e@��ti�?�            @l@�       �                   P`@r�q��?�             k@�       �       	             �?�t`�4 �?J            �^@������������������������       �                     �?�       �                    @8@W"�h�?I            @^@�       �                    �?��(\���?H             ^@�       �                   �W@������?	             .@������������������������       �                     @������������������������       �                     &@�       �                   i@���N8�??            @Z@������������������������       �                    �G@�       �                    �?��ϭ�*�?&             M@�       �                    �L@4��?�?#             J@�       �                   �_@؇���X�?            �A@�       �                   pp@�q�q�?             .@�       �                    �?����X�?             @������������������������       �                     �?�       �                   @]@r�q��?             @������������������������       �                     @�       �                    _@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     4@������������������������       �                     1@������������������������       �                     @������������������������       �                     �?�       �                    �?V��N��?<            �W@�       �                   �Z@F�t�K��?#            �L@�       �                   0a@      �?             @������������������������       �                     �?������������������������       �                     @�       �       	          033@f1r��g�?             �J@�       �       	          033@x�����?            �C@�       �                   p`@�MI8d�?            �B@������������������������       �                     �?�       �                   pb@4?,R��?             B@�       �                    �N@�t����?             A@�       �                     M@"pc�
�?             6@�       �       	          ����?      �?
             0@�       �                   �j@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                   @d@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     (@�       �                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        	             ,@�       �                   b@؀�:M�?            �B@�       �                    �H@r�q��?             @�       �                    a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       	             @¦	^_�?             ?@�       �                    X@�\��N��?             3@������������������������       �                      @�       �                    �L@��.k���?             1@�       �       	          ����?�<ݚ�?             "@�       �                     I@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �                   �`@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     (@�       �                   �X@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                    �M@,sI�v�?6            �V@�       �       	          ����?      �?             D@������������������������       �                     @�       �                    @J@�t����?             A@������������������������       �                     .@�       �       	          ����?�\��N��?             3@�       �                    @M@�<ݚ�?             "@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    �?�z�G��?	             $@�       �                    e@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�              	          ����?p���?             I@�       �                   �m@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                    �E@�t�bh�h(h+K ��h-��R�(KMKK��h^�B       �t@     �x@      o@     �]@      "@      H@       @     �@@              9@       @       @              @       @      @       @                      @      @      .@      �?      *@              "@      �?      @              @      �?      �?      �?                      �?      @       @      @                       @      n@     �Q@     �c@      :@     �E@      1@     �E@      .@       @       @       @       @       @      @              @       @      �?      �?              �?      �?              �?      �?                      @      @             �A@      @      A@      @      @      @      @      �?       @               @      �?      �?      �?              �?      �?              �?                       @      >@       @      @      �?      @      �?      @                      �?       @              8@      �?      4@              @      �?              �?      @              �?       @               @      �?                       @      ]@      "@      @      @      @                      @     @\@      @     �[@      @     �W@      �?      @@      �?      *@      �?      (@              �?      �?      �?                      �?      3@             �O@              .@       @      &@              @       @              �?      @      �?      @                      �?      @      @      @                      @     @T@     �F@      $@      <@      �?              "@      <@      �?      $@      �?      @      �?      @              @      �?                      �?              @       @      2@      @      @      @              @      @               @      @       @               @      @               @      ,@      �?      �?      �?                      �?      �?      *@      �?      @      �?       @               @      �?                       @              "@     �Q@      1@              @     �Q@      ,@      M@      @      @      @      @              �?      @      �?                      @     �I@       @     �I@      �?      E@              "@      �?      @               @      �?              �?       @                      �?      *@       @      *@      @      (@       @      @       @               @      @              "@              �?      �?              �?      �?                      @     �U@     �q@     �R@      i@      >@      4@      8@       @              @      8@      @      @      @      @                      @      4@              @      (@              (@      @             �F@     �f@      B@     �f@      &@     �[@      �?              $@     �[@      "@     �[@      @      &@      @                      &@      @      Y@             �G@      @     �J@      @     �G@      @      >@      @      $@      @       @              �?      @      �?      @               @      �?              �?       @                       @              4@              1@              @      �?              9@     @Q@      &@      G@      @      �?              �?      @               @     �F@       @      ?@      @      ?@      �?              @      ?@      @      >@      @      2@      �?      .@      �?      @              @      �?                      $@      @      @      @                      @              (@      �?      �?      �?                      �?       @                      ,@      ,@      7@      @      �?      �?      �?              �?      �?              @              "@      6@      "@      $@               @      "@       @      @       @      �?       @               @      �?              @               @      @              @       @      @       @                      @              (@      "@      �?              �?      "@              &@     �S@      $@      >@              @      $@      8@              .@      $@      "@      @       @      @      �?      @                      �?              �?      @      @      @      �?      @                      �?              @      �?     �H@      �?      @              @      �?                     �E@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK녔h}�Bh3         P                   P`@U�ք�?�           ��@       /                    �?j=M>�:�?�            �s@                           �?X�Emq�?A            �Z@                           `@r֛w���?             ?@������������������������       �                     "@                           �?���|���?
             6@������������������������       �                     @       	       	          ����?      �?             0@������������������������       �                     (@
                            P@      �?             @������������������������       �                      @������������������������       �                      @                          �\@�sly47�?/            �R@                          @X@8�Z$���?            �C@������������������������       �                     $@                           �E@V�a�� �?             =@������������������������       �                     @              	          ����?ȵHPS!�?             :@                          �Y@r�q��?             2@                           ]@      �?             @������������������������       �                      @                           �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@������������������������       �                      @       (                   `n@)O���?             B@       #       	          `ff�?��H�}�?             9@       "                    �H@���y4F�?             3@       !                    �?X�<ݚ�?             "@                            �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     $@$       '                    �?r�q��?             @%       &                    \@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @)       .                    �?�C��2(�?             &@*       -       	             �?�q�q�?             @+       ,                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @0       C                   P`@���ȑ��?             j@1       B                    �?ȵHPS!�?2            �S@2       5                    �?��ɉ�?*            @P@3       4       	             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?6       =                   `_@�8��8��?'             N@7       8                   (p@ ��WV�?!             J@������������������������       �                    �D@9       :                    @L@"pc�
�?             &@������������������������       �                      @;       <                    _@�q�q�?             @������������������������       �                     �?������������������������       �                      @>       ?                    �K@      �?              @������������������������       �                     @@       A                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@D       O                    �R@�z�N��?M            ``@E       F                   0q@ ����?L            @`@������������������������       �        <             Y@G       J                    �G@��S�ۿ?             >@H       I       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?K       N       	             �?h�����?             <@L       M                   �b@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     8@������������������������       �                     �?Q       �       	          ��� @@<QR���?           0z@R       �                    �?*2��`B�?�            Px@S       `                    �D@6�Nӆ�?a            �b@T       _                   �r@�LQ�1	�?             7@U       ^                   �f@�C��2(�?             6@V       W                   `]@���N8�?             5@������������������������       �                     &@X       ]                   �l@ףp=
�?             $@Y       Z                   �[@      �?             @������������������������       �                      @[       \                    a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?a       ~                    �?P�B�y��?P            @_@b       y                   �a@�LQ�1	�?+            @Q@c       v                   ``@�BbΊ�?&             M@d       e                   `T@#z�i��?            �D@������������������������       �                     @f       m                    �?      �?             B@g       h                    �?���Q��?             .@������������������������       �                     @i       j                   `\@���Q��?             $@������������������������       �                     @k       l                   @f@�q�q�?             @������������������������       �                      @������������������������       �                     @n       u                   �s@؇���X�?             5@o       t                    `P@ףp=
�?             4@p       s                   �k@�}�+r��?             3@q       r                   pj@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?������������������������       �                     �?w       x                   �x@�IєX�?             1@������������������������       �        
             0@������������������������       �                     �?z       {                   pb@"pc�
�?             &@������������������������       �                     @|       }                    �L@�q�q�?             @������������������������       �                      @������������������������       �                     @       �                    �?Dc}h��?%             L@�       �                   `a@v�2t5�?            �D@�       �                   �b@�ՙ/�?             5@�       �                   �g@��.k���?             1@�       �                   @_@�����H�?             "@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     @�       �                    @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �s@z�G�z�?             4@�       �                   �b@�����H�?             2@�       �                    �?@4և���?
             ,@�       �                   �a@      �?             @�       �                   @m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     .@�       �                   h@�p�?�             n@�       �                    �?��t���?�            �m@�       �                    �?�7��?0            �S@�       �                    �?`����֜?+            �Q@������������������������       �        '             O@�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �                    b@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �d@��G�?e            �c@�       �                    �?��[�8��?b             c@�       �       	          ����?����Q8�?.            �Q@�       �                   �a@P����?&            �M@�       �                   �\@@4և���?             ,@������������������������       �                     �?������������������������       �                     *@������������������������       �                    �F@�       �                   l@      �?             (@������������������������       �                     @�       �       	          `ff�?      �?             @�       �                    �?      �?             @������������������������       �                     �?�       �                   xp@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    @H�U?B�?4            �T@�       �                   @[@���!pc�?&            �K@������������������������       �                     @�       �       	          `ff�?�θ�?%             J@�       �                   `a@Jm_!'1�?#            �H@������������������������       �        	             &@�       �                     H@�I�w�"�?             C@������������������������       �                     0@�       �                     N@8�A�0��?             6@�       �                   �b@     ��?             0@������������������������       �                     @�       �                   �l@�z�G��?             $@������������������������       �                     @�       �       	          ����?      �?             @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                     I@|��?���?             ;@�       �                   �l@ףp=
�?             $@�       �                   `f@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �p@�t����?	             1@�       �                   �`@$�q-�?             *@�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     @�       �                    a@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �h@      �?             @������������������������       �                     @������������������������       �                     �?�       �       	          033@ףp=
�?             >@������������������������       �        
             ,@�       �                    �G@     ��?             0@�       �                   (p@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?$�q-�?             *@������������������������       �                     &@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h^�B�        t@     �y@      M@     p@      G@      N@      7@       @      "@              ,@       @              @      ,@       @      (@               @       @               @       @              7@      J@      @     �@@              $@      @      7@      @              @      7@      @      .@      @      @       @              �?      @      �?                      @              (@               @      1@      3@      0@      "@      .@      @      @      @       @      @              @       @              @              $@              �?      @      �?      �?      �?                      �?              @      �?      $@      �?       @      �?      �?              �?      �?                      �?               @      (@     �h@      "@     @Q@      "@      L@      @      �?      @                      �?      @     �K@       @      I@             �D@       @      "@               @       @      �?              �?       @              @      @              @      @      �?      @                      �?              *@      @      `@       @      `@              Y@       @      <@      �?      �?      �?                      �?      �?      ;@      �?      @      �?                      @              8@      �?             �p@     `c@     Pp@      `@     @P@     �T@      @      4@       @      4@      �?      4@              &@      �?      "@      �?      @               @      �?      �?      �?                      �?              @      �?              �?              O@     �O@     �F@      8@     �E@      .@      ;@      ,@              @      ;@      "@      "@      @      @              @      @              @      @       @               @      @              2@      @      2@       @      2@      �?       @      �?       @                      �?      $@                      �?              �?      0@      �?      0@                      �?       @      "@              @       @      @       @                      @      1@     �C@      1@      8@      *@       @      "@       @       @      �?      @              �?      �?              �?      �?              �?      @              @      �?      �?      �?                      �?      @              @      0@       @      0@      �?      *@      �?      @      �?      �?              �?      �?                       @              $@      �?      @              @      �?               @                      .@     �h@     �F@     `h@      E@     �R@      @     @Q@      �?      O@              @      �?              �?      @              @      @      @              �?      @              @      �?             @^@      C@      ^@     �@@     �P@      @      M@      �?      *@      �?              �?      *@             �F@              "@      @      @              @      @      �?      @              �?      �?       @               @      �?               @             �J@      =@      D@      .@              @      D@      (@      D@      "@      &@              =@      "@      0@              *@      "@      @      "@              @      @      @      @              �?      @      �?      �?              �?      �?                       @      @                      @      *@      ,@      �?      "@      �?      @      �?                      @              @      (@      @      (@      �?       @      �?              �?       @              $@                      @      �?      @      �?                      @      �?      @              @      �?              @      ;@              ,@      @      *@       @      �?       @                      �?      �?      (@              &@      �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuMhvh(h+K ��h-��R�(KM��h}�B88         �                    �?0����?�           ��@       A                    �?���\�?�            �x@                          @_@�E��
��?\            �c@                           �?�{��?��?"             K@������������������������       �                      @                           �?D>�Q�?              J@                          �Q@$�q-�?            �C@������������������������       �                      @	                           V@�?�|�?            �B@
              	          ����?���N8�?             5@              	          ���ܿ��S�ۿ?             .@������������������������       �                     @                          �Z@�C��2(�?             &@������������������������       �                     "@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        	             0@                            P@��
ц��?             *@                           �?���Q��?	             $@                           @L@؇���X�?             @                          `Y@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @       >                   �b@Np�����?:            �Y@       =                    �?��
ц��?5            �V@       2                   �n@~�hP��?,            �R@        +                   �c@z�G�z�?             D@!       "                    �?�X����?             6@������������������������       �                      @#       *       	          @33�?      �?             4@$       )                   �g@r�q��?             2@%       (                   @_@և���X�?             @&       '                    b@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     &@������������������������       �                      @,       -       	             �?�X�<ݺ?             2@������������������������       �                     (@.       /                     I@r�q��?             @������������������������       �                     @0       1       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?3       <                   �r@      �?             A@4       7                    �?��+7��?             7@5       6                   Pp@�q�q�?             @������������������������       �                      @������������������������       �                     �?8       ;                   @b@z�G�z�?             4@9       :                     N@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     ,@������������������������       �                     &@������������������������       �        	             1@?       @                   �a@���!pc�?             &@������������������������       �                     @������������������������       �                      @B       �                    �N@�����H�?�            `n@C       f                    �?��y�S��?x             h@D       S                    �I@ףp=
�?^            �b@E       R                   �e@ZՏ�m|�?!            �H@F       G                   �Z@��E�B��?             �G@������������������������       �                      @H       K                    �?�:�^���?            �F@I       J       	          ����?      �?             @������������������������       �                      @������������������������       �                      @L       Q       	          `ff�?������?            �D@M       N                    @G@      �?              @������������������������       �                     @O       P                   �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �@@������������������������       �                      @T       U                    �?�L�L��?=            @Y@������������������������       �                    �A@V       a                   @m@��IF�E�?+            �P@W       `                   `l@     ��?             @@X       Y                    �?�r����?             >@������������������������       �                     �?Z       _                   �`@ܷ��?��?             =@[       \                   �^@�θ�?	             *@������������������������       �                      @]       ^                   �j@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     0@������������������������       �                      @b       c                    @M@г�wY;�?             A@������������������������       �                     ?@d       e                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?g       t                    @M@�%^�?            �E@h       s                    �?؇���X�?             <@i       p       	             @z�G�z�?             4@j       k                   �[@r�q��?             2@������������������������       �                      @l       o                   �X@      �?
             0@m       n                   @^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@q       r       	             @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @u       x                    �?��S���?             .@v       w                   �s@���Q��?             @������������������������       �                      @������������������������       �                     @y       |                    �M@      �?             $@z       {                    _@z�G�z�?             @������������������������       �                     �?������������������������       �                     @}       �                   �a@z�G�z�?             @~                          �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �R@p���?              I@������������������������       �                     H@�       �                    a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          pff�?V~b���?�            �t@�       �                    I@J�:�Ȣ�?�            �o@�       �                   `_@      �?             0@�       �                    �?ףp=
�?             $@�       �                    `R@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    a@r�q��?             @������������������������       �                     @�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @��w\ud�?�            �m@�       �                    ]@�Cc}h��?�             l@�       �                   �Z@ �o_��?             9@������������������������       �                     @�       �                   `l@b�2�tk�?             2@������������������������       �                     @�       �                    �?���|���?             &@������������������������       �                     �?�       �                    �?�z�G��?             $@������������������������       �                     @�       �                    �D@      �?             @������������������������       �                      @�       �                   @[@      �?             @������������������������       �                      @�       �                     J@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �? l����?}            �h@�       �                   �j@H�_�r�?n            `f@������������������������       �        '            �P@�       �                    �?4�0_���?G            @\@�       �                   �^@ >�֕�?A            @Z@������������������������       �                    �C@�       �                    �?�C��2(�?,            �P@�       �       	            �?�(\����?             D@������������������������       �                    �A@�       �                    _@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   @o@���B���?             :@�       �                     G@���Q��?             $@������������������������       �                     @�       �                     M@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   `a@      �?             0@������������������������       �                     $@�       �       	          @33�?r�q��?             @�       �                   �t@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   pb@      �?              @�       �                   �`@      �?             @������������������������       �                      @�       �                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �]@�z�G��?             4@������������������������       �                     @�       �                   �`@      �?             0@������������������������       �                      @�       �                   `a@      �?              @������������������������       �                     @�       �                   Pc@      �?             @������������������������       �                      @������������������������       �                      @�       �                    @N@      �?
             ,@�       �                    �?���|���?             &@������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	          ���@^�JB=�?<            @T@�       �                   �d@�9mf��?,            �O@�       �                    �?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@�       �                    �?��e�B��?%            �I@�       �                    �?#z�i��?            �D@�       �                    �?$�q-�?             *@������������������������       �                     @�       �                   `o@      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �b@���>4��?             <@�       �                    a@����X�?
             ,@�       �                    @X�<ݚ�?             "@�       �                   @m@z�G�z�?             @�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �\@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   0e@d}h���?	             ,@�       �                    �?�8��8��?             (@�       �                    p@r�q��?             @������������������������       �                     @�       �                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �I@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                    �?�����H�?             2@������������������������       �                     �?�       �                    �?�IєX�?             1@������������������������       �                     *@�       �                    �?      �?             @������������������������       �                     �?�                           �P@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�b�B�      h�h(h+K ��h-��R�(KMKK��h^�B        u@     �x@     �V@     Ps@     �O@     @W@      &@     �E@       @              "@     �E@      @      B@       @              �?      B@      �?      4@      �?      ,@              @      �?      $@              "@      �?      �?              �?      �?                      @              0@      @      @      @      @      @      �?       @      �?              �?       @              @                      @              @      J@      I@     �H@      E@     �H@      9@      @@       @      .@      @               @      .@      @      .@      @      @      @       @      @       @                      @       @              &@                       @      1@      �?      (@              @      �?      @              �?      �?              �?      �?              1@      1@      @      1@       @      �?       @                      �?      @      0@      @       @      @                       @              ,@      &@                      1@      @       @      @                       @      ;@      k@      :@     �d@      .@     �`@       @     �D@      @     �D@       @              @     �D@       @       @       @                       @       @     �C@       @      @              @       @      �?              �?       @                     �@@       @              @     �W@             �A@      @     �M@      @      :@      @      :@      �?              @      :@      @      $@               @      @       @      @                       @              0@       @              �?     �@@              ?@      �?       @               @      �?              &@      @@      @      8@      @      0@      @      .@       @              �?      .@      �?       @               @      �?                      *@      �?      �?      �?                      �?               @      @       @       @      @       @                      @      @      @      @      �?              �?      @              �?      @      �?      �?              �?      �?                      @      �?     �H@              H@      �?      �?      �?                      �?     �n@     @V@     �j@     �C@      @      $@      �?      "@      �?       @               @      �?                      @      @      �?      @              �?      �?      �?                      �?      j@      =@     @i@      6@      2@      @      @              &@      @      @              @      @      �?              @      @              @      @      @       @              �?      @               @      �?      �?              �?      �?              g@      .@     @e@      "@     �P@              Z@      "@     �X@      @     �C@              N@      @     �C@      �?     �A@              @      �?              �?      @              5@      @      @      @      @              �?      @              @      �?              .@      �?      $@              @      �?      @      �?      @                      �?       @              @      @      �?      @               @      �?      �?      �?                      �?      @              ,@      @              @      ,@       @       @              @       @      @               @       @               @       @              @      @      @      @      @                      @      @              ?@      I@      =@      A@      �?      &@      �?                      &@      <@      7@      ;@      ,@      (@      �?      @              @      �?      @               @      �?       @                      �?      .@      *@      @      $@      @      @      �?      @      �?      �?              �?      �?                      @      @      �?              �?      @                      @      &@      @      &@      �?      @      �?      @              �?      �?              �?      �?              @                       @      �?      "@      �?                      "@       @      0@      �?              �?      0@              *@      �?      @              �?      �?       @      �?                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KKᅔh}�B81         l                   �`@�+	G�?�           ��@       Y                    �?l�"�^%�?�            �u@       .       	          ����?0�	B��?�            �n@       )                   `_@D�n�3�?;            �W@                            J@��(@��?-            �Q@                           �?      �?             4@                          �^@X�<ݚ�?             "@������������������������       �                     @	                           @H@�q�q�?             @
                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     &@       "                   �k@��H�}�?!             I@                          `c@�s��:��?             C@                           �?��<b���?             7@������������������������       �                     *@                           �?      �?             $@                          �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?և���X�?             @                          �]@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @                           �L@z�G�z�?
             .@������������������������       �                     @       !                    @M@�q�q�?             "@                           @Z@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @#       $                    �?�8��8��?             (@������������������������       �                     "@%       (                   @_@�q�q�?             @&       '                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?*       -                    �?H%u��?             9@+       ,                   �]@�nkK�?             7@������������������������       �                     �?������������������������       �                     6@������������������������       �                      @/       8                    �?h�˹�?g             c@0       1                    i@�����?             3@������������������������       �                      @2       7                    @������?
             1@3       4                   �]@@4և���?             ,@������������������������       �                     &@5       6                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @9       L                    �?ՀJ��?[            �`@:       A                    @M@io8�?N             ]@;       <       	          033@�(�Tw�?3            �S@������������������������       �        +             Q@=       >                    �?ףp=
�?             $@������������������������       �                      @?       @                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?B       K                    �O@�S����?             C@C       H                   P`@����X�?             5@D       G       	          ����?      �?             0@E       F                    @O@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @I       J                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     1@M       N                     I@�t����?             1@������������������������       �                     @O       X                    @�n_Y�K�?
             *@P       W                    c@�q�q�?	             (@Q       R                   �o@���!pc�?             &@������������������������       �                     @S       T                   �q@���Q��?             @������������������������       �                      @U       V                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?Z       _                    �?�C��2(�?A            �X@[       \                   �b@�q�q�?             "@������������������������       �                     @]       ^                    �?      �?             @������������������������       �                     @������������������������       �                     �?`       a                   �k@��S�ۿ?<            �V@������������������������       �        '             L@b       c                    @G@@�0�!��?             A@������������������������       �                      @d       g                   pm@      �?             @@e       f                    �P@      �?             @������������������������       �                      @������������������������       �                      @h       i                   �S@@4և���?             <@������������������������       �                     �?j       k                    �R@ 7���B�?             ;@������������������������       �                     :@������������������������       �                     �?m       �                    �?�E���?�            @x@n       s                   @E@��ʫf_�?�            �r@o       p                    �N@���N8�?             5@������������������������       �                     3@q       r                    �?      �?              @������������������������       �                     �?������������������������       �                     �?t       �                    �?2L�����?�            @q@u       z                    �?��W3�?*            �Q@v       w                   �b@PN��T'�?             ;@������������������������       �                     6@x       y                   0d@z�G�z�?             @������������������������       �                     @������������������������       �                     �?{       �                    �L@d�
��?             F@|       �       	          ����?�LQ�1	�?             7@}       �                   �d@���!pc�?             &@~       �                    e@�����H�?             "@       �                     F@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     (@�       �                   �l@؇���X�?             5@�       �       	          033@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     0@�       �                   ht@6��m�?�            �i@�       �       	          `ff@�DÓ ��?�            @i@�       �                   �]@(l58��?            �h@�       �                   �a@��R[s�?            �A@������������������������       �                     @�       �                    f@�חF�P�?             ?@�       �                    �?�GN�z�?             6@������������������������       �                     "@�       �                   pd@�n_Y�K�?
             *@�       �                     D@z�G�z�?             $@������������������������       �                     �?�       �                   �n@�����H�?             "@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                    @������?h            �d@�       �                    �?`-�I�w�?a             c@�       �                    f@ �Cc}�?             <@�       �                     N@�8��8��?             8@�       �                   �_@���N8�?             5@�       �                   pk@r�q��?             @�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �        
             .@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �f@      �?             @������������������������       �                     �?������������������������       �                     @�       �       	            �?�&/�E�?O             _@�       �                    �?@��8��??             X@�       �                    �?��f�{��?8            �U@������������������������       �        2             S@�       �                    �G@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �       	          ����?ףp=
�?             $@�       �                   �b@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?�>4և��?             <@�       �                    _@��<b���?             7@�       �                   �^@���Q��?             @�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   �b@�����H�?	             2@�       �                   �f@�IєX�?             1@������������������������       �                     �?������������������������       �                     0@������������������������       �                     �?������������������������       �                     @�       �                   �`@      �?             (@������������������������       �                     @�       �                    �?      �?              @�       �                     P@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �b@�DC��,�?2            �V@�       �                   �\@ 	��p�?!             M@�       �                   �m@���Q��?             $@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     H@�       �       	          ����?4���C�?            �@@�       �                    �?�<ݚ�?	             2@������������������������       �                     $@�       �                   �p@      �?              @������������������������       �                     @������������������������       �                     @�       �                    �?�q�q�?             .@�       �                   �p@r�q��?             (@������������������������       �                     $@������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h^�B       `t@     �y@     �T@     �p@     @R@     �e@     �K@      D@     �@@     �B@      .@      @      @      @              @      @       @      �?       @      �?                       @      @              &@              2@      @@      1@      5@      @      2@              *@      @      @       @      �?              �?       @              @      @      @       @      @                       @               @      (@      @      @              @      @       @      @       @                      @      @              �?      &@              "@      �?       @      �?      �?      �?                      �?              �?      6@      @      6@      �?              �?      6@                       @      2@     �`@      @      *@       @              @      *@      �?      *@              &@      �?       @      �?                       @      @              (@     @^@      @     @[@      �?     @S@              Q@      �?      "@               @      �?      �?      �?                      �?      @      @@      @      .@       @      ,@       @      @              @       @                      @      @      �?              �?      @                      1@      @      (@              @      @       @      @       @      @       @              @      @       @       @              �?       @      �?                       @      �?              �?              "@     �V@      @      @              @      @      �?      @                      �?      @      U@              L@      @      <@       @              @      <@       @       @               @       @               @      :@      �?              �?      :@              :@      �?             �n@      b@     �k@      S@      �?      4@              3@      �?      �?              �?      �?             �k@      L@      G@      9@      7@      @      6@              �?      @              @      �?              7@      5@      4@      @       @      @       @      �?       @      �?              �?       @              @                       @      (@              @      2@      @       @      @                       @              0@     �e@      ?@     �e@      <@     �e@      9@      :@      "@              @      :@      @      1@      @      "@               @      @       @       @              �?       @      �?      @      �?      @                      �?      @                      @      "@             �b@      0@     �a@      $@      9@      @      6@       @      4@      �?      @      �?       @      �?       @                      �?      @              .@               @      �?       @                      �?      @      �?              �?      @             @]@      @     �W@       @     @U@      �?      S@              "@      �?              �?      "@              "@      �?      @      �?              �?      @              @              7@      @      2@      @       @      @       @      �?              �?       @                       @      0@       @      0@      �?              �?      0@                      �?      @              @      @      @               @      @      �?      @              @      �?              �?                      @              @      7@      Q@      @      K@      @      @      @      �?              �?      @                      @              H@      3@      ,@      ,@      @      $@              @      @      @                      @      @      $@       @      $@              $@       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK�h}�B(5         �                    �?6������?�           ��@                           �?(��3Ea�?�             w@                          �R@N1���?'            �N@������������������������       �                     "@                           �J@��
ц��?!             J@                          `c@z�G�z�?             9@              	          ����?r�q��?             8@������������������������       �        
             3@	       
                   �`@z�G�z�?             @������������������������       �                     @                          Pn@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                           �P@l��
I��?             ;@              	          ����?�㙢�c�?             7@              	          @33�?X�<ݚ�?             "@������������������������       �                     @                            P@�q�q�?             @                           �?z�G�z�?             @                           �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �        	             ,@������������������������       �                     @       [                    �?N��s�?�            0s@       N       	          ����?�{���2�?M            �[@       A                   ``@P��E��?/             R@       <                    �?�q����?#            �J@        ;                    @O@��]�T��?            �D@!       :                   �f@��Q��?             D@"       9                    �?�����?             C@#       8                   po@��R[s�?            �A@$       7                   �k@�q�q�?             ;@%       6       	             �? �o_��?             9@&       -                   `Z@�q�q�?             8@'       ,                   @E@և���X�?             @(       )                   �_@���Q��?             @������������������������       �                      @*       +                     L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @.       /                   �h@@�0�!��?             1@������������������������       �                     "@0       3                    �?      �?              @1       2                   Pa@      �?              @������������������������       �                     �?������������������������       �                     �?4       5                   �b@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?=       >                   �l@�8��8��?             (@������������������������       �                     "@?       @       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?B       K                    �?�����?             3@C       J       	             �?X�Cc�?             ,@D       E                     E@�q�q�?             (@������������������������       �                      @F       I                    m@�z�G��?             $@G       H                   �^@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @L       M                    @P@z�G�z�?             @������������������������       �                     @������������������������       �                     �?O       Z                   �t@�ݜ�?            �C@P       Y                    �?�L���?            �B@Q       R                   �U@؇���X�?             5@������������������������       �                      @S       X                    @K@�}�+r��?             3@T       U                    �J@�����H�?             "@������������������������       �                     @V       W                   �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@������������������������       �                     0@������������������������       �                      @\       �                   �d@Hm_!'1�?�            �h@]       �                    �R@�v�|�<�?            �g@^       _                   �U@8v�YeK�?~            �g@������������������������       �                      @`       �                   0c@��ɹ?}            �g@a       �                   0c@x��-�?j            �c@b       �                   Hq@Х-��ٹ?d            �b@c       d                    �F@T(y2��?O            �]@������������������������       �                     6@e       p       	          hff�?DE�SA_�?B            @X@f       o                   �b@      �?             0@g       h                   �_@؇���X�?             ,@������������������������       �                      @i       n                   �^@�q�q�?             @j       k                    �O@z�G�z�?             @������������������������       �                     @l       m                   0o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @q       z                   @l@H�!b	�?6            @T@r       s                    �M@ pƵHP�?#             J@������������������������       �                    �@@t       u       	          ����?�}�+r��?             3@������������������������       �                     &@v       y       	             @      �?              @w       x                   @`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @{       �                    �?ܷ��?��?             =@|                           @G@ �Cc}�?             <@}       ~       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `\@$�q-�?             :@�       �                   `[@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �        
             0@������������������������       �                     �?������������������������       �                     ?@�       �                   �p@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     =@������������������������       �                     �?�       �                   Pe@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?H��Ly��?�            �v@�       �       	          ���@��11��?�            �r@�       �                   Hp@T;���?�            �q@�       �                   �c@�P�U`��?�            `h@�       �       	          ����?�G��l��?             5@�       �                    @���!pc�?             &@�       �                   �_@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �_@z�G�z�?             $@�       �                   `^@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?�8���?y            �e@������������������������       �        <            @T@�       �                    Z@��a�n`�?=            @W@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @L@����\�?:            �V@�       �                   Pd@      �?,             P@������������������������       �                     A@�       �                   �n@��S�ۿ?             >@�       �                   m@h�����?             <@������������������������       �                     6@�       �                   @m@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?���B���?             :@�       �                    d@      �?             8@�       �                   �l@�IєX�?	             1@������������������������       �                     &@�       �                   �l@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �       	          033�?����X�?             @�       �                   �i@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �?Z��:���?1            �V@�       �       	          ����?HP�s��?             9@������������������������       �                     3@�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?8�A�0��?             �P@�       �                   �d@�-ῃ�?            �N@�       �                    d@�����?            �L@�       �       	          ����?�xGZ���?            �A@�       �                    @��X��?             <@�       �                   Pa@�㙢�c�?             7@������������������������       �                     $@�       �       	          ����?�	j*D�?             *@�       �                   �c@���Q��?             $@�       �                    �K@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   `]@�C��2(�?             6@������������������������       �                      @������������������������       �                     4@������������������������       �                     @������������������������       �                     @�       �                   �i@$�q-�?	             *@������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �b@P�~D&�?+            �P@�       �                   �r@PN��T'�?#             K@�       �                    �J@�8��8��?             H@�       �                    �?�θ�?             *@������������������������       �                      @�       �                    `@�C��2(�?             &@������������������������       �                      @�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	          ����?��?^�k�?            �A@�       �                    _@@4և���?             ,@������������������������       �                     &@�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     5@�       �                   �a@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �C@�θ�?             *@������������������������       �                     @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK�KK��h^�B0       �t@     �x@     �S@      r@      <@     �@@              "@      <@      8@      4@      @      4@      @      3@              �?      @              @      �?      �?      �?                      �?              �?       @      3@      @      3@      @      @              @      @       @      @      �?      �?      �?              �?      �?              @                      �?              ,@      @              I@     p@      A@     @S@      =@     �E@      0@     �B@      .@      :@      ,@      :@      (@      :@      "@      :@      "@      2@      @      2@      @      1@      @      @       @      @               @       @      �?       @                      �?       @              @      ,@              "@      @      @      �?      �?      �?                      �?       @      @              @       @                      �?       @                       @      @               @              �?              �?      &@              "@      �?       @               @      �?              *@      @      "@      @      @      @               @      @      @      @      @              @      @              @               @              @      �?      @                      �?      @      A@      @      A@      @      2@       @              �?      2@      �?       @              @      �?       @               @      �?                      $@              0@       @              0@     �f@      *@     @f@      (@     @f@       @              $@     @f@      $@     �b@       @     �a@       @     �[@              6@       @     @V@      @      (@       @      (@               @       @      @      �?      @              @      �?      �?              �?      �?              �?               @              @     @S@      �?     �I@             �@@      �?      2@              &@      �?      @      �?      @      �?                      @              @      @      :@      @      9@      �?      �?      �?                      �?       @      8@       @       @               @       @                      0@              �?              ?@       @      @              @       @                      =@      �?              @       @      @                       @     p@     @[@     �m@      N@     �m@      H@      f@      3@      &@      $@      @       @      @       @               @      @                      @       @       @       @       @       @                       @      @             �d@      "@     @T@              U@      "@      �?       @      �?                       @     �T@      @      O@       @      A@              <@       @      ;@      �?      6@              @      �?              �?      @              �?      �?              �?      �?              5@      @      5@      @      0@      �?      &@              @      �?              �?      @              @       @       @       @               @       @              @                       @      O@      =@      7@       @      3@              @       @               @      @             �C@      ;@     �C@      6@     �C@      2@      3@      0@      3@      "@      3@      @      $@              "@      @      @      @      �?      @      �?                      @      @              @                      @              @      4@       @               @      4@                      @              @      �?      (@               @      �?      @      �?                      @      2@     �H@       @      G@      @      F@      @      $@       @              �?      $@               @      �?       @      �?                       @      �?      A@      �?      *@              &@      �?       @      �?                       @              5@      @       @      @                       @      $@      @              @      $@        �t�bubhhubehhub.